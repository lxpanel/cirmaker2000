CircuitMaker Text
5.6
Probes: 1
v2[p]
Operating Point
0 180 227 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 40 30 100 10
197 87 1865 1000
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.499458 0.500000
365 183 478 280
9437202 0
0
6 Title:
5 Name:
0
0
0
22
13 Logic Switch~
5 647 600 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
45097.7 1
0
13 Logic Switch~
5 644 682 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
45097.7 0
0
13 Logic Switch~
5 372 360 0 1 11
0 14
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V11
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
45097.7 3
0
13 Logic Switch~
5 375 278 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V10
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3421 0 0
2
45097.7 2
0
14 Logic Display~
6 1082 682 0 1 2
10 2
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 L8
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8157 0 0
2
45097.7 0
0
10 2-In NAND~
219 1022 686 0 3 22
0 4 3 2
0
0 0 624 0
4 7400
-7 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
5572 0 0
2
45097.7 0
0
14 Logic Display~
6 1080 642 0 1 2
10 5
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 L5
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8901 0 0
2
45097.7 0
0
8 2-In OR~
219 904 649 0 3 22
0 3 4 5
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U2A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
7361 0 0
2
45097.7 0
0
9 2-In NOR~
219 740 614 0 3 22
0 7 4 3
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U1B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
4747 0 0
2
45097.7 5
0
9 2-In NOR~
219 741 692 0 3 22
0 3 6 4
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U1A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
972 0 0
2
45097.7 4
0
14 Logic Display~
6 896 612 0 1 2
10 3
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 L4
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3472 0 0
2
45097.7 3
0
14 Logic Display~
6 893 699 0 1 2
21 4
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 L3
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9998 0 0
2
45097.7 2
0
12 Hex Display~
7 416 179 0 18 19
10 15 14 13 12 0 0 0 0 0
0 1 1 1 1 0 1 1 9
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
3536 0 0
2
45097.7 13
0
14 Logic Display~
6 621 377 0 1 2
21 12
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 L7
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4597 0 0
2
45097.7 12
0
14 Logic Display~
6 624 290 0 1 2
10 13
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 L6
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3835 0 0
2
45097.7 11
0
9 2-In NOR~
219 469 370 0 3 22
0 13 14 12
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U4B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
3670 0 0
2
45097.7 10
0
9 2-In NOR~
219 468 292 0 3 22
0 15 12 13
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
5616 0 0
2
45097.7 9
0
9 2-In NOR~
219 935 297 0 3 22
0 11 8 9
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U4C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
9323 0 0
2
45097.7 8
0
9 2-In NOR~
219 936 375 0 3 22
0 9 10 8
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U4D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
317 0 0
2
45097.7 7
0
14 Logic Display~
6 1091 295 0 1 2
10 9
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 L1
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3108 0 0
2
45097.7 6
0
14 Logic Display~
6 1088 382 0 1 2
21 8
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 L2
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4299 0 0
2
45097.7 5
0
8 Hex Key~
166 883 185 0 11 12
0 11 10 9 8 0 0 0 0 0
1 49
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
9672 0 0
2
45097.7 4
0
30
1 3 2 0 0 8320 0 5 6 0 0 4
1066 686
1046 686
1046 686
1049 686
0 2 3 0 0 8320 0 0 6 8 0 5
872 616
872 689
990 689
990 695
998 695
0 1 4 0 0 4224 0 0 6 5 0 4
870 678
885 678
885 677
998 677
1 3 5 0 0 4224 0 7 8 0 0 4
1064 646
948 646
948 649
937 649
0 2 4 0 0 0 0 0 8 7 0 3
870 703
870 658
891 658
0 1 3 0 0 0 0 0 8 8 0 3
865 616
865 640
891 640
0 1 4 0 0 0 0 0 12 12 0 4
791 692
841 692
841 703
877 703
0 1 3 0 0 0 0 0 11 11 0 3
811 614
811 616
880 616
1 2 6 0 0 12416 0 2 10 0 0 4
656 682
688 682
688 701
728 701
1 1 7 0 0 4224 0 1 9 0 0 4
659 600
721 600
721 605
727 605
3 1 3 0 0 128 0 9 10 0 0 6
779 614
811 614
811 718
720 718
720 683
728 683
3 2 4 0 0 128 0 10 9 0 0 6
780 692
791 692
791 647
710 647
710 623
727 623
4 0 8 0 0 8320 0 22 0 0 17 4
874 209
874 355
1028 355
1028 375
3 0 9 0 0 8320 0 22 0 0 18 4
880 209
880 277
1046 277
1046 299
2 2 10 0 0 4224 0 22 19 0 0 7
886 209
886 349
877 349
877 370
910 370
910 384
923 384
1 1 11 0 0 4224 0 22 18 0 0 7
892 209
892 268
891 268
891 283
914 283
914 288
922 288
0 1 8 0 0 0 0 0 21 20 0 4
986 375
1036 375
1036 386
1072 386
0 1 9 0 0 0 0 0 20 19 0 3
1006 297
1006 299
1075 299
3 1 9 0 0 0 0 18 19 0 0 6
974 297
1006 297
1006 401
915 401
915 366
923 366
3 2 8 0 0 0 0 19 18 0 0 6
975 375
986 375
986 330
905 330
905 306
922 306
4 0 12 0 0 8320 0 13 0 0 25 4
407 203
407 350
561 350
561 370
3 0 13 0 0 8320 0 13 0 0 26 4
413 203
413 272
579 272
579 294
2 0 14 0 0 4224 0 13 0 0 27 4
419 203
419 344
405 344
405 360
1 0 15 0 0 4096 0 13 0 0 28 4
425 203
425 263
424 263
424 278
0 1 12 0 0 0 0 0 14 30 0 4
519 370
569 370
569 381
605 381
0 1 13 0 0 0 0 0 15 29 0 3
539 292
539 294
608 294
1 2 14 0 0 0 0 3 16 0 0 4
384 360
416 360
416 379
456 379
1 1 15 0 0 4224 0 4 17 0 0 4
387 278
449 278
449 283
455 283
3 1 13 0 0 0 0 17 16 0 0 6
507 292
539 292
539 396
448 396
448 361
456 361
3 2 12 0 0 0 0 16 17 0 0 6
508 370
519 370
519 325
438 325
438 301
455 301
17
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
1102 689 1219 713
1112 697 1208 713
12 inverse stat
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
1097 616 1214 640
1107 624 1203 640
12 primary stat
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
589 669 634 693
599 677 623 693
3 SET
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
571 585 632 609
581 593 621 609
5 RESET
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
890 570 967 594
900 578 956 594
7 primary
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
894 709 971 733
904 717 960 733
7 inverse
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
630 37 811 61
640 45 800 61
20 Set-Reset (SR) Latch
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 17
641 56 798 80
651 64 787 80
17 (its like memory)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
1084 162 1185 186
1094 170 1174 186
10 state here
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 19
921 162 1094 186
931 170 1083 186
19 <<-- type in memory
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
964 97 1089 121
974 105 1078 121
13 3 = no memory
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
619 330 696 354
629 338 685 354
7 inverse
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
618 248 695 272
628 256 684 272
7 primary
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
299 263 360 287
309 271 349 287
5 RESET
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
317 347 362 371
327 355 351 371
3 SET
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
1085 253 1162 277
1095 261 1151 277
7 primary
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
1086 335 1163 359
1096 343 1152 359
7 inverse
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
