CircuitMaker Text
5.6
Probes: 1
v2[p]
Operating Point
0 180 227 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
209 87 1877 1000
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.499458 0.500000
377 183 490 280
9437202 0
0
6 Title:
5 Name:
0
0
0
37
13 Logic Switch~
5 921 494 0 1 11
0 15
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V11
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3965 0 0
2
45097.4 0
0
13 Logic Switch~
5 924 412 0 10 11
0 16 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V10
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8239 0 0
2
45097.4 1
0
13 Logic Switch~
5 228 474 0 1 11
0 23
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
828 0 0
2
45097.4 2
0
13 Logic Switch~
5 224 387 0 1 11
0 19
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6187 0 0
2
45097.4 3
0
13 Logic Switch~
5 230 322 0 1 11
0 24
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7107 0 0
2
45097.4 4
0
13 Logic Switch~
5 1100 284 0 1 11
0 26
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6433 0 0
2
45097.4 5
0
13 Logic Switch~
5 1096 217 0 1 11
0 27
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8559 0 0
2
45097.4 6
0
13 Logic Switch~
5 705 200 0 1 11
0 29
0
0 0 21360 0
2 0V
-8 13 6 21
2 V4
-6 24 8 32
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3674 0 0
2
5.90082e-315 0
0
13 Logic Switch~
5 665 183 0 1 11
0 30
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5697 0 0
2
5.90082e-315 5.26354e-315
0
13 Logic Switch~
5 189 226 0 1 11
0 31
0
0 0 21360 0
2 0V
-6 -18 8 -10
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3805 0 0
2
5.90082e-315 5.30499e-315
0
13 Logic Switch~
5 197 186 0 1 11
0 32
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5219 0 0
2
5.90082e-315 5.32571e-315
0
9 2-In AND~
219 698 778 0 3 22
0 12 11 10
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
3795 0 0
2
45097.5 0
0
10 Ascii Key~
169 653 639 0 11 12
0 12 9 8 7 6 5 4 3 0
1 49
0
0 0 4656 0
0
4 KBD2
-14 -34 14 -26
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 0 0 0 0 0
3 KBD
3637 0 0
2
45097.5 0
0
10 Ascii Key~
169 557 641 0 11 12
0 11 34 35 36 37 38 39 40 0
0 49
0
0 0 4656 0
0
4 KBD1
-14 -34 14 -26
0
0
0
0
0
4 SIP8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
0 0 0 512 0 0 0 0
3 KBD
3226 0 0
2
45097.5 0
0
14 Ascii Display~
172 855 713 0 42 44
0 4 5 6 7 8 9 10 3 0
28 12849 12849 12850 12336 12336 12593 12593 12336 12336
12336 12336 12337 12593 12593 8224 8224 8224 8224 8224
8224 8224 8224 8224 8224 8224 8224 8224 8224 8224
8224 8224 8224
0
0 0 21104 0
4 1MEG
-15 -42 13 -34
5 DISP1
-3 -48 32 -40
0
0
102 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
%DE %5 0 %V
%DF %6 0 %V
%DG %7 0 %V
%DH %8 0 %V
0
0
0
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
82 0 0 0 0 0 0 0
4 DISP
6966 0 0
2
45097.4 0
0
14 Logic Display~
6 1170 511 0 1 2
10 13
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 L7
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9796 0 0
2
45097.4 0
0
14 Logic Display~
6 1173 424 0 1 2
10 14
0
0 0 53872 270
6 100MEG
3 -16 45 -8
2 L6
-5 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5952 0 0
2
45097.4 0
0
9 2-In NOR~
219 1018 504 0 3 22
0 14 15 13
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U4B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
3649 0 0
2
45097.4 9
0
9 2-In NOR~
219 1017 426 0 3 22
0 16 13 14
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3716 0 0
2
45097.4 10
0
7 Ground~
168 732 497 0 1 3
0 2
0
0 0 53360 90
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4797 0 0
2
45097.4 11
0
7 Ground~
168 662 345 0 1 3
0 2
0
0 0 53360 90
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4681 0 0
2
45097.4 12
0
5 4030~
219 506 344 0 3 22
0 22 23 18
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U3C
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 3 0
1 U
9730 0 0
2
45097.4 13
0
5 4030~
219 373 335 0 3 22
0 24 19 22
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U3B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 3 0
1 U
9874 0 0
2
45097.4 14
0
8 2-In OR~
219 575 498 0 3 22
0 21 20 17
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U2B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
364 0 0
2
45097.4 15
0
9 2-In AND~
219 446 452 0 3 22
0 22 23 21
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
3656 0 0
2
45097.4 16
0
9 2-In AND~
219 384 502 0 3 22
0 24 19 20
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
3131 0 0
2
45097.4 17
0
7 Ground~
168 1389 235 0 1 3
0 2
0
0 0 53360 90
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6772 0 0
2
45097.4 18
0
5 4030~
219 1208 240 0 3 22
0 27 26 25
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U3A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 3 0
1 U
9557 0 0
2
45097.4 19
0
7 Ground~
168 967 189 0 1 3
0 2
0
0 0 53360 90
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5789 0 0
2
5.90082e-315 5.34643e-315
0
8 2-In OR~
219 825 191 0 3 22
0 30 29 28
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U2A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
7328 0 0
2
5.90082e-315 5.3568e-315
0
7 Ground~
168 516 206 0 1 3
0 2
0
0 0 53360 90
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4799 0 0
2
5.90082e-315 5.36716e-315
0
9 2-In AND~
219 357 207 0 3 22
0 32 31 33
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
9196 0 0
2
5.90082e-315 5.37752e-315
0
5 Lamp~
206 665 488 0 2 3
11 17 2
0
0 0 624 0
3 100
-10 -24 11 -16
2 L5
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
3857 0 0
2
45097.4 22
0
5 Lamp~
206 585 334 0 2 3
11 18 2
0
0 0 624 0
3 100
-10 -24 11 -16
2 L4
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
7125 0 0
2
45097.4 23
0
5 Lamp~
206 1320 224 0 2 3
11 25 2
0
0 0 624 0
3 100
-10 -24 11 -16
2 L3
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
3641 0 0
2
45097.4 24
0
5 Lamp~
206 910 178 0 2 3
11 28 2
0
0 0 624 0
3 100
-10 -24 11 -16
2 L2
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
9821 0 0
2
5.90082e-315 5.38788e-315
0
5 Lamp~
206 456 194 0 2 3
11 33 2
0
0 0 624 0
3 100
-10 -24 11 -16
2 L1
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 L
3187 0 0
2
5.90082e-315 5.39306e-315
0
43
8 0 3 0 0 12416 0 13 0 0 11 6
632 663
631 663
631 732
708 732
708 742
719 742
7 1 4 0 0 8320 0 13 15 0 0 3
638 663
638 682
789 682
6 2 5 0 0 8320 0 13 15 0 0 3
644 663
644 691
789 691
5 3 6 0 0 8320 0 13 15 0 0 3
650 663
650 700
789 700
4 4 7 0 0 8320 0 13 15 0 0 3
656 663
656 709
789 709
3 5 8 0 0 8320 0 13 15 0 0 3
662 663
662 718
789 718
2 6 9 0 0 8320 0 13 15 0 0 3
668 663
668 727
789 727
3 7 10 0 0 4224 0 12 15 0 0 4
719 778
773 778
773 736
789 736
1 2 11 0 0 4224 0 14 12 0 0 3
578 665
578 787
674 787
1 1 12 0 0 4224 0 13 12 0 0 2
674 663
674 769
0 8 3 0 0 128 0 0 15 0 0 4
716 742
731 742
731 744
783 744
0 1 13 0 0 4096 0 0 16 17 0 4
1068 504
1118 504
1118 515
1154 515
0 1 14 0 0 8192 0 0 17 16 0 3
1088 426
1088 428
1157 428
1 2 15 0 0 12416 0 1 18 0 0 4
933 494
965 494
965 513
1005 513
1 1 16 0 0 4224 0 2 19 0 0 4
936 412
998 412
998 417
1004 417
3 1 14 0 0 8320 0 19 18 0 0 6
1056 426
1088 426
1088 530
997 530
997 495
1005 495
3 2 13 0 0 12416 0 18 19 0 0 6
1057 504
1068 504
1068 459
987 459
987 435
1004 435
2 1 2 0 0 4096 0 33 20 0 0 3
677 501
725 501
725 498
2 1 2 0 0 8320 0 34 21 0 0 3
597 347
597 346
655 346
3 1 17 0 0 8320 0 24 33 0 0 3
608 498
608 501
653 501
3 1 18 0 0 8320 0 22 34 0 0 3
539 344
539 347
573 347
1 0 19 0 0 8192 0 4 0 0 23 3
236 387
236 388
321 388
2 2 19 0 0 8320 0 23 26 0 0 4
357 344
321 344
321 511
360 511
3 2 20 0 0 4224 0 26 24 0 0 4
405 502
547 502
547 507
562 507
3 1 21 0 0 4224 0 25 24 0 0 4
467 452
528 452
528 489
562 489
0 1 22 0 0 4224 0 0 25 27 0 3
409 335
409 443
422 443
3 1 22 0 0 0 0 23 22 0 0 2
406 335
490 335
0 2 23 0 0 4096 0 0 25 29 0 2
404 461
422 461
2 1 23 0 0 12416 0 22 3 0 0 4
490 353
404 353
404 474
240 474
0 1 24 0 0 4224 0 0 26 31 0 3
337 326
337 493
360 493
1 1 24 0 0 0 0 5 23 0 0 4
242 322
265 322
265 326
357 326
1 2 2 0 0 0 0 27 35 0 0 3
1382 236
1382 237
1332 237
3 1 25 0 0 4224 0 28 35 0 0 4
1241 240
1296 240
1296 237
1308 237
1 2 26 0 0 4224 0 6 28 0 0 4
1112 284
1182 284
1182 249
1192 249
1 1 27 0 0 4224 0 7 28 0 0 4
1108 217
1184 217
1184 231
1192 231
2 1 2 0 0 0 0 36 29 0 0 3
922 191
960 191
960 190
3 1 28 0 0 4224 0 30 36 0 0 2
858 191
898 191
1 2 29 0 0 4224 0 8 30 0 0 2
717 200
812 200
1 1 30 0 0 4224 0 9 30 0 0 3
677 183
812 183
812 182
1 2 31 0 0 4224 0 10 32 0 0 4
201 226
325 226
325 216
333 216
1 1 32 0 0 4224 0 11 32 0 0 4
209 186
318 186
318 198
333 198
1 2 2 0 0 0 0 31 37 0 0 2
509 207
468 207
3 1 33 0 0 4224 0 32 37 0 0 2
378 207
444 207
12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
983 332 1164 356
993 340 1153 356
20 Set-Reset (SR) Latch
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
866 481 911 505
876 489 900 505
3 SET
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
848 397 909 421
858 405 898 421
5 RESET
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
404 265 505 289
414 273 494 289
10 Full Adder
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
739 483 800 507
749 491 789 507
5 CARRY
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
672 331 717 355
682 339 706 355
3 SUM
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
1135 106 1220 130
1145 114 1209 130
8 xor gate
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
301 107 386 131
311 115 375 131
8 and gate
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
779 96 856 120
789 104 845 120
7 or gate
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
1167 382 1244 406
1177 390 1233 406
7 primary
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
1168 464 1245 488
1178 472 1234 488
7 inverse
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 17
1097 559 1254 583
1107 567 1243 583
17 (its like memory)
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
